module Control(
    Op_i       ,
    ID_EX_o,
    PC_i_mux_o,
    branch_o
);
input[5:0]      Op_i;
output[7:0]     ID_EX_o;
output          PC_i_mux_o;
output          branch_o;


endmodule
